LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_arith.ALL;
USE IEEE.STD_LOGIC_unsigned.ALL;
USE IEEE.numeric_std.ALL;

ENTITY UART_TXHEAD_EN_BLOCK IS

    PORT (
        i_Addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        i_BaseAddr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        o_En : OUT STD_LOGIC := '0'
    );
END UART_TXHEAD_EN_BLOCK;

ARCHITECTURE arch OF UART_TXHEAD_EN_BLOCK IS

    CONSTANT UART0 : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0000";
    CONSTANT UART1 : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0800";
    CONSTANT UART2 : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"1000";
    CONSTANT UART3 : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"1800";
    CONSTANT UART4 : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"2000";
    CONSTANT UART5 : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"2800";

    CONSTANT RXDATA : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0000";
    CONSTANT TXDATA : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0200";
    CONSTANT RXTAIL : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0400";
    CONSTANT RXHEAD : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0401";
    CONSTANT TXTAIL : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0402";
    CONSTANT TXHEAD : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0403";
    CONSTANT CTRL : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0408";

BEGIN

    o_En <= '1' WHEN (i_Addr = i_BaseAddr + TXHEAD) ELSE
        '0';

END arch;