-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 9.1 Build 350 03/24/2010 Service Pack 2 SJ Web Edition"
-- CREATED		"Thu Jul 04 14:44:46 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY one_wire_module IS 
	PORT
	(
		DATA_WR_READY :  IN  STD_LOGIC;
		MHz_25 :  IN  STD_LOGIC;
		DATA_RE_READY :  IN  STD_LOGIC;
		OW_IN :  IN  STD_LOGIC;
		kHz :  IN  STD_LOGIC;
		MHz :  IN  STD_LOGIC;
		BASE_ADDR :  IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		DATA_FROM_MPU :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		MPU_ADDR :  IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		OW_OUT :  OUT  STD_LOGIC;
		DATA_TO_MPU :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END one_wire_module;

ARCHITECTURE bdf_type OF one_wire_module IS 

COMPONENT dpram_1wire_name
	PORT(wren : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 rdaddress : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 wraddress : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dpram_1wire_temp
	PORT(wren : IN STD_LOGIC;
		 rden : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 rdaddress : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 wraddress : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT tri31_1
	PORT(enabledt : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 tridata : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT one_wire_block_v3
	PORT(i_Clk : IN STD_LOGIC;
		 i_MHz : IN STD_LOGIC;
		 i_kHz : IN STD_LOGIC;
		 i_1WIRE : IN STD_LOGIC;
		 i_DataRD : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 o_WR : OUT STD_LOGIC;
		 o_1WIRE : OUT STD_LOGIC;
		 o_AddrRD : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 o_AddrWR : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 o_DataWR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_Test : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	ADDR_EN :  STD_LOGIC;
SIGNAL	ADDR_RD_NAME :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	DATA_TO_MPU_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(63 DOWNTO 0);


BEGIN 



b2v_inst : dpram_1wire_name
PORT MAP(wren => SYNTHESIZED_WIRE_0,
		 clock => SYNTHESIZED_WIRE_1,
		 data => DATA_FROM_MPU,
		 rdaddress => ADDR_RD_NAME,
		 wraddress => MPU_ADDR(4 DOWNTO 0),
		 q => SYNTHESIZED_WIRE_22);


SYNTHESIZED_WIRE_2 <= NOT(MPU_ADDR(14) XOR BASE_ADDR(14));


SYNTHESIZED_WIRE_8 <= NOT(MPU_ADDR(8) XOR BASE_ADDR(8));


SYNTHESIZED_WIRE_11 <= NOT(MPU_ADDR(5) XOR BASE_ADDR(5));


SYNTHESIZED_WIRE_5 <= NOT(MPU_ADDR(11) XOR BASE_ADDR(11));


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_2 AND SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_4 AND SYNTHESIZED_WIRE_5;


SYNTHESIZED_WIRE_9 <= NOT(MPU_ADDR(7) XOR BASE_ADDR(7));


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_6 AND SYNTHESIZED_WIRE_7 AND SYNTHESIZED_WIRE_8 AND SYNTHESIZED_WIRE_9;


SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_10 AND SYNTHESIZED_WIRE_11;


SYNTHESIZED_WIRE_23 <= DATA_RE_READY AND ADDR_EN;


SYNTHESIZED_WIRE_6 <= NOT(MPU_ADDR(10) XOR BASE_ADDR(10));


b2v_inst24 : dpram_1wire_temp
PORT MAP(wren => SYNTHESIZED_WIRE_12,
		 rden => SYNTHESIZED_WIRE_23,
		 clock => SYNTHESIZED_WIRE_14,
		 data => SYNTHESIZED_WIRE_15,
		 rdaddress => MPU_ADDR(3 DOWNTO 0),
		 wraddress => SYNTHESIZED_WIRE_16,
		 q => SYNTHESIZED_WIRE_18);


b2v_inst26 : tri31_1
PORT MAP(enabledt => SYNTHESIZED_WIRE_23,
		 data => SYNTHESIZED_WIRE_18,
		 tridata => DATA_TO_MPU_ALTERA_SYNTHESIZED);


SYNTHESIZED_WIRE_10 <= NOT(MPU_ADDR(6) XOR BASE_ADDR(6));


ADDR_EN <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_0 <= DATA_WR_READY AND ADDR_EN;


SYNTHESIZED_WIRE_1 <= NOT(MHz_25);



SYNTHESIZED_WIRE_14 <= NOT(MHz_25);



b2v_inst6 : one_wire_block_v3
PORT MAP(i_Clk => MHz_25,
		 i_MHz => MHz,
		 i_kHz => kHz,
		 i_1WIRE => OW_IN,
		 i_DataRD => SYNTHESIZED_WIRE_22,
		 o_WR => SYNTHESIZED_WIRE_12,
		 o_1WIRE => OW_OUT,
		 o_AddrRD => ADDR_RD_NAME,
		 o_AddrWR => SYNTHESIZED_WIRE_16,
		 o_DataWR => SYNTHESIZED_WIRE_15);


SYNTHESIZED_WIRE_3 <= NOT(MPU_ADDR(13) XOR BASE_ADDR(13));


SYNTHESIZED_WIRE_4 <= NOT(MPU_ADDR(12) XOR BASE_ADDR(12));


SYNTHESIZED_WIRE_7 <= NOT(MPU_ADDR(9) XOR BASE_ADDR(9));

DATA_TO_MPU <= DATA_TO_MPU_ALTERA_SYNTHESIZED;

END bdf_type;