-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 9.1 Build 350 03/24/2010 Service Pack 2 SJ Web Edition"
-- CREATED		"Thu Jul 04 14:46:50 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY uart_module IS 
	PORT
	(
		RO_REZ :  IN  STD_LOGIC;
		RO_OSN :  IN  STD_LOGIC;
		DATA_WR_READY :  IN  STD_LOGIC;
		MHz_25 :  IN  STD_LOGIC;
		DATA_RE_READY :  IN  STD_LOGIC;
		BASE_ADDR :  IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		DATA_FROM_MPU :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		DQMBn :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		MPU_ADDR :  IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		DI_OSN :  OUT  STD_LOGIC;
		DI_REZ :  OUT  STD_LOGIC;
		NRE :  OUT  STD_LOGIC;
		DATA_TO_MPU :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		TEST :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END uart_module;

ARCHITECTURE bdf_type OF uart_module IS 

COMPONENT uart_rxhead_en_block
	PORT(i_Addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_BaseAddr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 o_En : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT uart_txhead_block
	PORT(i_Clk : IN STD_LOGIC;
		 i_En : IN STD_LOGIC;
		 i_Addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_BaseAddr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_Data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_TxHead : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uart_txtail_en_block
	PORT(i_Addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_BaseAddr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 o_En : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT uart_txdata_block
	PORT(i_Clk : IN STD_LOGIC;
		 i_TxStart : IN STD_LOGIC;
		 i_DriverReady : IN STD_LOGIC;
		 i_MPU_RE : IN STD_LOGIC;
		 i_DataReadyWE : IN STD_LOGIC;
		 i_Addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_MPU_Data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 i_RamData : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 i_TxHead : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 o_RamRE : OUT STD_LOGIC;
		 o_DV : OUT STD_LOGIC;
		 o_RamAddr : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		 o_TxData : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 o_TxTail : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uart_rx_block
	PORT(i_Clk : IN STD_LOGIC;
		 i_Rx : IN STD_LOGIC;
		 o_RxDV : OUT STD_LOGIC;
		 o_RxData : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uart_rxdata_block
	PORT(i_Clk : IN STD_LOGIC;
		 i_DV : IN STD_LOGIC;
		 i_DataReadyWE : IN STD_LOGIC;
		 i_MPU_Data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 i_RxData : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 o_RamWE : OUT STD_LOGIC;
		 o_ByteSel : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 o_RamAddr : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		 o_RamData : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_RxHead : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dpram_2k
	PORT(wren : IN STD_LOGIC;
		 rden : IN STD_LOGIC;
		 inclock : IN STD_LOGIC;
		 outclock : IN STD_LOGIC;
		 byteena_a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 rdaddress : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 wraddress : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT tri31_1
	PORT(enabledt : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 tridata : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uart_ctrl_block
	PORT(i_Clk : IN STD_LOGIC;
		 i_En : IN STD_LOGIC;
		 i_Addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_BaseAddr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_Data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_Mode : OUT STD_LOGIC;
		 o_Loopback : OUT STD_LOGIC;
		 o_Channel : OUT STD_LOGIC;
		 o_TxStart : OUT STD_LOGIC;
		 o_CtrlReg : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uart_txhead_en_block
	PORT(i_Addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_BaseAddr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 o_En : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT uart_ctrl_en_block
	PORT(i_Addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 i_BaseAddr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 o_En : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT uart_tx_block
	PORT(i_Clk : IN STD_LOGIC;
		 i_TxDV : IN STD_LOGIC;
		 i_Data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 o_TX : OUT STD_LOGIC;
		 o_TX_Active : OUT STD_LOGIC;
		 o_Ready : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT mux1
	PORT(data1 : IN STD_LOGIC;
		 data0 : IN STD_LOGIC;
		 sel : IN STD_LOGIC;
		 result : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	ByteSel_WR :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	CHANNEL :  STD_LOGIC;
SIGNAL	CLK :  STD_LOGIC;
SIGNAL	CTRL :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	DATA_EN :  STD_LOGIC;
SIGNAL	DATA_TO_MPU_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	DI :  STD_LOGIC;
SIGNAL	DI_OSN_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	DI_REZ_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	DRIVER_READY :  STD_LOGIC;
SIGNAL	LOOPBACK :  STD_LOGIC;
SIGNAL	MODE :  STD_LOGIC;
SIGNAL	NRE_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	RAM_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	RAM_RD_ADDR :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	RAM_RE :  STD_LOGIC;
SIGNAL	RAM_TO_MPU_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	RAM_WE :  STD_LOGIC;
SIGNAL	RAM_WR_ADDR :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	RAM_WR_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	RX_DATA :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	RX_DV :  STD_LOGIC;
SIGNAL	RX_HEAD :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	RXHEAD_ADDR_EN :  STD_LOGIC;
SIGNAL	TEST_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	TX_DATA :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	TX_DV :  STD_LOGIC;
SIGNAL	TX_TAIL :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	TX_WE :  STD_LOGIC;
SIGNAL	TXHEAD :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	TXSTART :  STD_LOGIC;
SIGNAL	TXTAIL_ADDR_EN :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_0 <= NOT(MPU_ADDR(14) XOR BASE_ADDR(14));


b2v_inst11 : uart_rxhead_en_block
PORT MAP(i_Addr => MPU_ADDR,
		 i_BaseAddr => BASE_ADDR,
		 o_En => RXHEAD_ADDR_EN);


SYNTHESIZED_WIRE_3 <= NOT(MPU_ADDR(11) XOR BASE_ADDR(11));


DATA_EN <= SYNTHESIZED_WIRE_0 AND SYNTHESIZED_WIRE_1 AND SYNTHESIZED_WIRE_2 AND SYNTHESIZED_WIRE_3;


b2v_inst14 : uart_txhead_block
PORT MAP(i_Clk => MHz_25,
		 i_En => DATA_WR_READY,
		 i_Addr => MPU_ADDR,
		 i_BaseAddr => BASE_ADDR,
		 i_Data => DATA_FROM_MPU,
		 o_TxHead => TXHEAD);


b2v_inst15 : uart_txtail_en_block
PORT MAP(i_Addr => MPU_ADDR,
		 i_BaseAddr => BASE_ADDR,
		 o_En => TXTAIL_ADDR_EN);


b2v_inst16 : uart_txdata_block
PORT MAP(i_Clk => CLK,
		 i_TxStart => TXSTART,
		 i_DriverReady => DRIVER_READY,
		 i_MPU_RE => DATA_RE_READY,
		 i_DataReadyWE => SYNTHESIZED_WIRE_4,
		 i_Addr => MPU_ADDR,
		 i_MPU_Data => DATA_FROM_MPU,
		 i_RamData => RAM_DATA,
		 i_TxHead => TXHEAD(10 DOWNTO 0),
		 o_RamRE => RAM_RE,
		 o_DV => TX_DV,
		 o_RamAddr => RAM_RD_ADDR,
		 o_TxData => TX_DATA,
		 o_TxTail => TX_TAIL);


SYNTHESIZED_WIRE_23 <= DATA_RE_READY AND DATA_EN AND SYNTHESIZED_WIRE_5;

TEST_ALTERA_SYNTHESIZED(0) <= CLK;


TEST_ALTERA_SYNTHESIZED(1) <= DI_OSN_ALTERA_SYNTHESIZED;


TEST_ALTERA_SYNTHESIZED(2) <= DI_REZ_ALTERA_SYNTHESIZED;


TEST_ALTERA_SYNTHESIZED(3) <= RO_OSN;



b2v_inst22 : uart_rx_block
PORT MAP(i_Clk => CLK,
		 i_Rx => SYNTHESIZED_WIRE_6,
		 o_RxDV => RX_DV,
		 o_RxData => RX_DATA);


b2v_inst23 : uart_rxdata_block
PORT MAP(i_Clk => CLK,
		 i_DV => RX_DV,
		 i_DataReadyWE => SYNTHESIZED_WIRE_7,
		 i_MPU_Data => DATA_FROM_MPU,
		 i_RxData => RX_DATA,
		 o_RamWE => RAM_WE,
		 o_ByteSel => ByteSel_WR,
		 o_RamAddr => RAM_WR_ADDR,
		 o_RamData => RAM_WR_DATA,
		 o_RxHead => RX_HEAD);

TEST_ALTERA_SYNTHESIZED(4) <= RO_REZ;



b2v_inst25 : dpram_2k
PORT MAP(wren => RAM_WE,
		 rden => SYNTHESIZED_WIRE_23,
		 inclock => SYNTHESIZED_WIRE_24,
		 outclock => SYNTHESIZED_WIRE_24,
		 byteena_a => ByteSel_WR,
		 data => RAM_WR_DATA,
		 rdaddress => MPU_ADDR(8 DOWNTO 0),
		 wraddress => RAM_WR_ADDR,
		 q => RAM_TO_MPU_DATA);


b2v_inst26 : tri31_1
PORT MAP(enabledt => SYNTHESIZED_WIRE_11,
		 data => RX_HEAD,
		 tridata => DATA_TO_MPU_ALTERA_SYNTHESIZED);


b2v_inst27 : tri31_1
PORT MAP(enabledt => SYNTHESIZED_WIRE_12,
		 data => RAM_TO_MPU_DATA,
		 tridata => DATA_TO_MPU_ALTERA_SYNTHESIZED);


b2v_inst28 : tri31_1
PORT MAP(enabledt => SYNTHESIZED_WIRE_13,
		 data => TX_TAIL,
		 tridata => DATA_TO_MPU_ALTERA_SYNTHESIZED);


b2v_inst29 : dpram_2k
PORT MAP(wren => TX_WE,
		 rden => RAM_RE,
		 inclock => SYNTHESIZED_WIRE_25,
		 outclock => SYNTHESIZED_WIRE_25,
		 byteena_a => DQMBn,
		 data => DATA_FROM_MPU,
		 rdaddress => RAM_RD_ADDR,
		 wraddress => MPU_ADDR(8 DOWNTO 0),
		 q => RAM_DATA);


b2v_inst3 : uart_ctrl_block
PORT MAP(i_Clk => MHz_25,
		 i_En => DATA_WR_READY,
		 i_Addr => MPU_ADDR,
		 i_BaseAddr => BASE_ADDR,
		 i_Data => DATA_FROM_MPU,
		 o_Mode => MODE,
		 o_Channel => CHANNEL,
		 o_TxStart => TXSTART,
		 o_CtrlReg => CTRL);

TEST_ALTERA_SYNTHESIZED(5) <= NRE_ALTERA_SYNTHESIZED;


TEST_ALTERA_SYNTHESIZED(6) <= RX_DATA(1);


TEST_ALTERA_SYNTHESIZED(7) <= RX_DATA(0);



b2v_inst33 : uart_txhead_en_block
PORT MAP(i_Addr => MPU_ADDR,
		 i_BaseAddr => BASE_ADDR,
		 o_En => SYNTHESIZED_WIRE_16);


b2v_inst34 : tri31_1
PORT MAP(enabledt => SYNTHESIZED_WIRE_16,
		 data => TXHEAD,
		 tridata => DATA_TO_MPU_ALTERA_SYNTHESIZED);


b2v_inst35 : uart_ctrl_en_block
PORT MAP(i_Addr => MPU_ADDR,
		 i_BaseAddr => BASE_ADDR,
		 o_En => SYNTHESIZED_WIRE_17);


b2v_inst36 : tri31_1
PORT MAP(enabledt => SYNTHESIZED_WIRE_17,
		 data => CTRL,
		 tridata => DATA_TO_MPU_ALTERA_SYNTHESIZED);


SYNTHESIZED_WIRE_20 <= NOT(MPU_ADDR(10) OR SYNTHESIZED_WIRE_18);


SYNTHESIZED_WIRE_5 <= NOT(MPU_ADDR(10) OR MPU_ADDR(9));


TX_WE <= DATA_WR_READY AND SYNTHESIZED_WIRE_19;


b2v_inst5 : uart_tx_block
PORT MAP(i_Clk => CLK,
		 i_TxDV => TX_DV,
		 i_Data => TX_DATA,
		 o_TX => DI,
		 o_TX_Active => NRE_ALTERA_SYNTHESIZED,
		 o_Ready => DRIVER_READY);


SYNTHESIZED_WIRE_19 <= DATA_EN AND SYNTHESIZED_WIRE_20;


DI_OSN_ALTERA_SYNTHESIZED <= DI OR CHANNEL;


SYNTHESIZED_WIRE_12 <= DATA_RE_READY AND SYNTHESIZED_WIRE_23;


CLK <= MODE AND MHz_25;


SYNTHESIZED_WIRE_25 <= NOT(MHz_25);



SYNTHESIZED_WIRE_13 <= DATA_RE_READY AND TXTAIL_ADDR_EN;


SYNTHESIZED_WIRE_4 <= DATA_WR_READY AND TXTAIL_ADDR_EN;


SYNTHESIZED_WIRE_18 <= NOT(MPU_ADDR(9));



SYNTHESIZED_WIRE_24 <= NOT(MHz_25);



SYNTHESIZED_WIRE_7 <= DATA_WR_READY AND RXHEAD_ADDR_EN;


SYNTHESIZED_WIRE_11 <= DATA_RE_READY AND RXHEAD_ADDR_EN;


DI_REZ_ALTERA_SYNTHESIZED <= DI OR SYNTHESIZED_WIRE_22;


SYNTHESIZED_WIRE_22 <= NOT(CHANNEL);



SYNTHESIZED_WIRE_1 <= NOT(MPU_ADDR(13) XOR BASE_ADDR(13));


SYNTHESIZED_WIRE_2 <= NOT(MPU_ADDR(12) XOR BASE_ADDR(12));


b2v_inst9 : mux1
PORT MAP(data1 => RO_REZ,
		 data0 => RO_OSN,
		 sel => CHANNEL,
		 result => SYNTHESIZED_WIRE_6);

DI_OSN <= DI_OSN_ALTERA_SYNTHESIZED;
DI_REZ <= DI_REZ_ALTERA_SYNTHESIZED;
NRE <= NRE_ALTERA_SYNTHESIZED;
DATA_TO_MPU <= DATA_TO_MPU_ALTERA_SYNTHESIZED;
TEST <= TEST_ALTERA_SYNTHESIZED;

END bdf_type;